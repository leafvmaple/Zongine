       P��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ''''''''''''''            '''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                            '''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                            ''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                            '''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                        '''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                    '''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                  ''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                ''''''''''''''''''''''''''''''''''''''''                                                                                                                  ''''''''                                                                                                                                                                                                                                                                                                              ''''''''''''''''''''''''''''''''''''''''                                                                                    '''''''''          '''''''''                                                                                                                                                                                                                                                                                                              '''''''''''''''''''''''''''''''''''''''''                                                                                '''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                            ''''''''''''''''''''''''''''''''''''''''''                                                                              '''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                            '''''''''''''''''''''''''''''''''''''''''''                                                                          ''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                            '''''''''''''''''''''''''''''''''''''''''''        '''''                                                        ''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                              ''''''''''''''''''''''''''''''''''''''''''  ''''''''                                                        '''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                          '''''''''''''''''''''''''''''''''''''''''''  ''''''''                                                        ''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                        '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                    ''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                    '''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                            '''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                              '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                        '''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                            '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''  '''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                          ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                        ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                              ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                        ''''''''''                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                    ''''''''''''                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                  ''''''''''''''                                                                                                                                                                                                                                    ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                ''''''''''''''                                                                                                                                                                                                                                      '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                          '''''''''''''''                                                                                                                                                                                                                                        '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                        '''''''''''''''                                                                                                                                                                                                                                        '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                  ''''''''''''''''                                                                                                                                                                                                                                            '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                              ''''''''''''''''                                                                                                                                                                                                                                              ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''            '''''''''''''''''''''                                                                                                                                                                                                                                                ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''          '''''''''''''''''''''                                                                                                                                                                                                                                                  ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''      ''''''''''''''''''''''                                                                                                                                                                                                                                                    ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                    '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                        ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                          '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                            ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                    ''''''''''''''''''''''''''''''  ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                        ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                        ''''''''''''''''''''''''''''''''''''''''''  '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                        ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                          ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                            ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                              '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                      '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                        '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                            ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                  ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                    ''''''''''''''''''''''''''''''''''''''''''''''''''  ''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                      ''''''''''''''''''''''''''''''''''''  '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                          ''''''''''''''''''''''''''''''''''    ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                              ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                      ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                            '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                    '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                          ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                            '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''  '''''''                                                                                                                                                                                                                                                                                                                                                                              '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                      '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                          '''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                        '''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                          ''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                      '''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                          '''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                              ''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                '''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                        ''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                      '''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                    '''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                      '''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                      '''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                            ''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                            ''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                ''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                ''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                        '''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                              '''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                          '''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                    '''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                      '''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                        ''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                          '''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                          '''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                              '''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                        ''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                              '''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                              '''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                      '''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                              '''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                ''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''              '''''''''                                                                              ''''''''                                                                                                                                                                                                                                                                                '''''''''''''''''''''''''''''''''''''''''''''''''''''''''          '''''''''''''''                                                                      ''''''''                                                                                                                                                                                                                                                                                '''''''''''''''''''''''''''''''''''''''''''''''''''''''''  '''''''''''''''''''''                                                                  ''''''''                                                                                                                                                                                                                                                                                          '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                            ''''''''                                                                                                                                                                                                                                                                                          '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                        ''''''''                                                                                                                                                                                                                                                                                                  ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                  ''''''''                                                                                                                                                                                                                                                                                                      ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                              ''''''''                                                                                                                                                                                                                                                                                                        '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                              ''''''''                                                                                                                                                                                                                                                                                                        ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                ''    ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                            ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                ''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                  '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                      '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                              '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                      '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                      ''''''''''''''''''''''''''''''''''''''              ''''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                      ''''''''''''''''''''''''''''''''''''''                  ''''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                      ''''''''''''''''''''''''''''''''''                            '''''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                      '''''''''''''''''''''''''''''''                                      '''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                      '''''''''''''''''''''''''''''''                                          '''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                            ''''''''''''''''''''''''''''                                      '''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                '''''''''''''''''''''''''''                                    '''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                  ''''''''''''''''''''''''''                                    '''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                    '''''''''''''''''''''''                                        '''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                  ''''''''''''''''''''''''                                        '''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                  ''''''''''''''''''''''''                                        '''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                  ''''''''''''''''''''''''                                        '''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                  ''''''''''''''''''''''''                                          ''''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                  ''''''''''''''''''''''                                                  ''''''''''''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''''''                                                        ''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                        ''''''''''''''''''                                                              '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                '''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            '''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      '''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  '''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        '''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      '''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      '''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ''''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          '''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ''''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            '''''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          '''''''''''''''''''                                                                                                                                  